
module D0_Pixel(MINUS, PLUS);
inout MINUS, PLUS;
endmodule
