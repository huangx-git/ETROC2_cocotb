
module ETROC2_Peripheral_Caps(
    VDD_QInj,
    VDD_PA,
    VDD_Dis,
    VDD_D,
    VDD_SL,
    VDD_CLK,
    VSS_QInj,
    VSS_PA,
    VSS_Dis,
    VSS_D,
    VSS_SL,
    VSS_CLK
);
inout VDD_QInj, VDD_PA, VDD_Dis, VDD_D, VDD_SL, VDD_CLK, VSS_QInj, VSS_PA, VSS_Dis, VSS_D, VSS_SL, VSS_CLK;

endmodule