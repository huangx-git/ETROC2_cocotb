
module D1_Pixel(MINUS, PLUS);
inout MINUS, PLUS;
endmodule
