
module DSUP(vss_IO, vdd_IO, vss, vdd);
inout vss_IO, vdd_IO, vss, vdd;


endmodule
