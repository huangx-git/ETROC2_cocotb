
module D2_Pixel(MINUS, PLUS);
inout MINUS, PLUS;
endmodule
