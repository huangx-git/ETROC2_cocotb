`timescale 1ns/1ps
module IOPWR(vss_IO, vdd_IO, vss);
inout vss_IO, vdd_IO, vss;
endmodule
