//Verilog HDL for "ETROC_PLL_Core_feedbackDivider", "majorityVoterBalanced"
//"functional"


module majorityVoterBalanced ( inA, inB, inC, out, tmrErr, VDD, VSS );


  parameter WIDTH = 1;
  input   [(WIDTH-1):0]   inA, inB, inC;
  output  [(WIDTH-1):0]   out;
  output                  tmrErr;
  inout VDD, VSS;
  reg                     tmrErr;
  assign out = (inA&inB) | (inA&inC) | (inB&inC);
  always @(inA or inB or inC)
  begin
    if (inA!=inB || inA!=inC || inB!=inC)
      tmrErr = 1;
    else
      tmrErr = 0;
  end

endmodule

