
module PixelCaps(
    VDD_QInj,
    VDD_PA,
    VDD_Dis,
    VDD_D,
    VSS_QInj,
    VSS_PA,
    VSS_Dis,
    VSS_D
);
inout     VDD_QInj,    VDD_PA,    VDD_Dis,     VDD_D,     VSS_QInj,     VSS_PA,     VSS_Dis,     VSS_D;

endmodule