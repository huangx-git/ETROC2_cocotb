../verification/CERN_IO_PAD_H_ECON.sv