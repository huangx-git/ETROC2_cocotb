
module D3_Pixel(MINUS, PLUS);
inout MINUS, PLUS;
endmodule
